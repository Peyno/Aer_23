package Tb; 

interface AufzugIfc; 

endinterface 


module mkAufzug(AufzugIfc); 

endmodule

endpackage