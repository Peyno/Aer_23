package Settings;
  Integer width = 1173;
  Integer height = 470;

  // Settings for graytest.png. Comment out the above settings and comment in the below ones.
  //Integer width = 16;
  //Integer height = 16;
  Integer n_vals = width * height;
endpackage