package AcceleratorChecker;
    import MyTypes::*;
    import GetPut::*;
    import ClientServer::*;
    import FIFO::*;
    import ImageFunctions::*;
    import Gauss::*;
    import StmtFSM::*;
    import Settings::*;
    import Vector::*;
    import GaussTop::*;
        

    module mkAcceleratorChecker(Empty);
        // TODO: implement me with a StmtFSM
    endmodule : mkAcceleratorChecker
endpackage : AcceleratorChecker